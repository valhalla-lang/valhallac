f : Int -> Int
f n = n - 20

a = 2 + f 3 * 4 / 6

-- Treat `3` literal as intger numeric in type checker.
