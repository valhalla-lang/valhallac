A <> B
(<>) A B
((<>) A) B

--      CALL
--      /  \
--     /    \
--   CALL    B
--   /  \
--  /    \
-- <>     A