!infix (+++) 20 :left
!posfix ~ 70

a = 3 +++ 2
b = a + 7~
