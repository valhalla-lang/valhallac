2 + 3.2  -- 2 natural gets cast to 2.0 real.
-3 + 4   -- 4 natural gets cased to 4 integer.
4 + 5    -- 4 and 5 stay natural.
