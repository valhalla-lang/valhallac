f : Int -> Int
f n = n - 20

a = 2 + f -3 * 4 / 6
