import :IO

IO::puts "Hello, World."
