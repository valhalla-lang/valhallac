subset I Int

(n, m) : I^2
