
ys = [| 2; 2; 3 |]

assert (ys == [| 2; 2; 3 |]
