[ :puts, print
  :gets, input ] = import :IO

name = input "> "
puts "Hello, " + name.captialise + "."

