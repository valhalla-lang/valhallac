a : Nat
a = 3

__raw_print (a + 2.5)

