a : Nat -> Nat -> Int
a n m = n - 2*m

a 1 2

-- a = n |-> (m |-> n - 2*m)
--           |_____________|
--                  |
--               func: `__a_final`
--     |_____________________|
--                |
--             func: `__a__0`
-- |__________________________|
--          |
--       func: a