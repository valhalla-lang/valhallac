3 + 4 * 2 - 1
-1 * 2

