a : Nat
a = 3  -- only one byte

__raw_print (a + 2.5)
__raw_print "hello"
