-- Without using the prelude, or importing IO...

_write_stream :1 "Hello, World.\n"
