f : A -> B -> C
a = n + 3