a : Nat
a = 0xabc

__raw_print (a + 2.5)

