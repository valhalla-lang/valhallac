a : Nat -> Nat -> Int
a n m = n - 2*m

a 1 2

-- a = n |-> (m |-> n - 2*m)
--           |_____________|
--                  |
--               func: `a__1`
--     |_____________________|
--                |
--             func: `a__0`
-- |__________________________|
--          |
--       func: a