a - b - c - d