a : Nat -> Nat -> Int
a n m = n + 2*m

a 1 2