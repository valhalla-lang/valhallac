2 + 3
-- same as
(+) 2 3
-- same as
(2 +) 3
-- same as
(+ 3) 2