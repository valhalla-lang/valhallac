2
34
2.3
-2