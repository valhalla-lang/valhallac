# Without using the prelude, or importing IO...

_write_stream :STDOUT "Hello, World.\n"
