a : Set Nat
a = Nat

b : a
b = 6 * 7