3 + 8 * 9