4 + 3
5 - 4
3 * 4.0
3 + :a
