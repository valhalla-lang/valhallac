a : Nat
a = 3 + 9

b : Real
b = a + 4

