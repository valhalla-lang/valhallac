(- a)
(+ a)
(* a)
