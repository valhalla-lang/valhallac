2 + 3.0   -- Constant folds to 5.0 (Real).

-4 + (10 + 2)  -- Folds to 8 (Natural).

3 + -2.0  -- Folds to 1.0 (Real).

(-) 2 3  -- Folds to -1 (Integer).

2 + 3 * 3 - 8 / 2.0   -- 7.0 (Real).