-2 3
