3 + 2; 1 - 89; 2 - 3 * 4
3 + 1
