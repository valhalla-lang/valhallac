(2 + 3)  -- Eq. of: ((2 +) 3), can write: ((+ 3) 2)
(2 +)
(+ 3)  -- Partial application


----
2 + 3
-- same as
(+) 2 3
-- same as
(2 +) 3
-- same as
(+ 3) 2