a : Int
a = 3 + 9