a = 3 + 6
b = a + 2