-- I is subset of the integers.
I <: Int
I : Power(Int) -- the same as above

-- n and m are both integers.
(n, m) : I^2
(n, m) : I*I  -- the same as above
