(2 + 3)  -- Eq. of: ((2 +) 3), can write: ((+ 3) 2)
(2 +)
(+ 3)  -- Partial application