n : Nat => n mod 3 is 0