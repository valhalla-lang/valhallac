a : Nat
a = 3 + 9

b : Real
b = a + 4

c : XyZ
c = hello (3 * 8)