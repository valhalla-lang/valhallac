- 8