f = 2
x = 4

x

f x