漢字 = "hello漢字漢字 world"
 漢字漢字   漢字v